----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:29:53 04/11/2013 
-- Design Name: 
-- Module Name:    UART - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity UART is
    Port ( clk : in  STD_LOGIC;
			  reset : in STD_LOGIC;
			  send : in STD_LOGIC;
           uart_input : in  STD_LOGIC_VECTOR (7 downto 0):="00000000";
           uart_output : out  STD_LOGIC_VECTOR (7 downto 0):="00000000");
			  
end UART;

architecture Behavioral of UART is

component Transmitter is
    Port ( input : in  STD_LOGIC_VECTOR (7 downto 0); --  the parallel input to transmitter module
           output : out  STD_LOGIC; 						-- the serial output generated by the transmitter module
           clk_in : in  STD_LOGIC; 							-- input clock to transmitter
           send : in  STD_LOGIC; 							-- send bit to load and start transfer of parallel input
           data_sent : out  STD_LOGIC; 					-- this is high when the 8 bits appended to low start bit are transmitted
           reset : in  STD_LOGIC); 							-- to reset the transmitter
end component;

component receiver is
    Port ( serial_input : in  STD_LOGIC; 						-- serial input to the receiver.
           clk : in  STD_LOGIC; 									-- Clock
			  reset :in  STD_LOGIC; 							-- reset the receiver to idle state
           output : out  STD_LOGIC_VECTOR (7 downto 0)); -- parallel output (8 bits) from the receiver.
			  
end component;



signal transmitted_output : std_logic :='1';
signal data_sent : std_logic :='0';
signal clk_192, clk_3072 : std_logic := '0';
signal count1, count2 : integer :=0;
begin


-- Map transmitter to UART module
tx : Transmitter 
Port Map ( 
	input => uart_input,						-- input to transmitter 
	output => transmitted_output,			-- transmitter output is stored temporarily
	clk_in => clk_192,						-- give 19.2 kHz clock as clock input
	send => send,								-- send bit to indicate when data received is to be given as output
	data_sent => data_sent,					-- data_sent is 1 when all data is transmitted
	reset => reset								-- reset is mapped to master reset 
);

-- Map receiver to UART module
rx : Receiver
Port Map (
	serial_input => transmitted_output,	-- take input from generated output
	clk => clk_3072,							-- 307.2 kHz clock
	reset => reset,							-- reset the receiver
	output => uart_output					-- output of UART
);

process(clk,clk_3072)
begin 

	-- when rising edge of clock, count till 162
	-- if count is 162 then reset the count
	 if (rising_edge(clk)) then
		if (count1 = 162) then 
			count1<=0;
			if (clk_3072 ='1') then
			clk_3072 <= '0';
			elsif (clk_3072 ='0') then
			clk_3072 <= '1';
			end if;
		else
			count1<=count1+1;
		end if;
	end if;

	-- when rising edge of clk_3072, count till 8
	-- if count is 8 then reset the count
		 if (rising_edge(clk_3072)) then
		if (count2 = 7) then 
			count2<=0;
			if (clk_192 ='1') then
			clk_192 <= '0';
			elsif (clk_192 ='0') then
			clk_192 <= '1';
			end if;
		else
			count2<=count2+1;
		end if;
	end if;
	
	


end process;



--count1 : Counter
--Generic Map (overflow_count => 163)
--Port Map (
--	reset => reset,
--	counter_clk => clk,
--	overflow => overflow1
--);
--
--count2 : Counter
--Generic Map (overflow_count => 8)
--Port Map (
--	reset => reset,
--	counter_clk => clk_3072,
--	overflow => overflow2
--);
--
--
--process(overflow1, overflow2)
--begin
--	if (overflow1'event) then 
--		if (clk_3072 ='1') then
--			clk_3072 <= '0';
--		elsif (clk_3072 ='0') then
--			clk_3072 <= '1';
--		end if;
--		report "Astha" severity note;
--	end if;
--	
--	if (overflow2='1') then
--		if (clk_192 ='1') then
--			clk_192 <= '0';
--		elsif (clk_192 ='0') then
--			clk_192 <= '1';
--		end if;
--		
--	end if;

-- end process;
	
end Behavioral;

