----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:33:07 04/11/2013 
-- Design Name: 
-- Module Name:    Transmitter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Transmitter is
    Port ( input : in  STD_LOGIC_VECTOR (7 downto 0); --  the parallel input to transmitter module
           output : out  STD_LOGIC; 						-- the serial output generated by the transmitter module
           clk_in : in  STD_LOGIC; 							-- input clock to transmitter
           send : in  STD_LOGIC; 							-- send bit to load and start transfer of parallel input
           data_sent : out  STD_LOGIC; 					-- this is high when the 8 bits appended to low start bit are transmitted
           reset : in  STD_LOGIC); 							-- to reset the transmitter
end Transmitter;

architecture Behavioral of Transmitter is

	 -- declaration of the PISO shifft register
	 COMPONENT PISO_shift_reg
    PORT(
         clk_s : IN  std_logic; 										-- input clock to PISO
         load : IN  std_logic; 										-- load input of PISO
         parallel_input : IN  std_logic_vector(7 downto 0); -- Parallel input to PISO
         serial_output : OUT  std_logic 							-- Serial output from PISO
        );
    END COMPONENT;
	 
	 -- declaration of Counter
	 COMPONENT Counter
	 Generic ( overflow_count : integer :=15 						-- default overflow count
				);
    PORT(
         reset : IN  std_logic; 										-- Counter reset 
         counter_clk : IN  std_logic; 								-- Clock to counter
         overflow : OUT  std_logic 									-- Overflow bit of counter
        );
    END COMPONENT;
    
-- States of transmitter:
-- Idle : when no output/input action is being performed
-- Start_transmission : Appending 0 bit to input when send is '1' (load the parallel input in register)
-- Data_transmission : Transmitting the 8 data bits (using counter and PISO)
-- Stop_transmission : Adding high bit to indicate completion of data transfer
type state is (idle, start_transmission, data_transmission, stop_transmission);
signal p_state, n_state : state :=idle; -- present and next state

signal load : std_logic := '0'; 				-- signal to load input to PISO
signal out_temp :std_logic := '1'; 			-- store the output of PISO to out_temp
signal overflow : std_logic := '0'; 		-- overflow bit to indicate overflow of counter (count till 8)
signal reset_counter : std_logic := '0'; 	-- reset the counter to 0


begin
	-- Port map of PISO shift register
	piso: PISO_shift_reg
	Port Map (
		clk_s => clk_in, 							-- the input clock is same as transmitter clock
      load => load, 								-- load input from transmitter signals
      parallel_input => input, 				-- input of PISO is given from input of transmitter
      serial_output => out_temp 				-- the output of PISO is stored to out_temp
	);
	
	--  
	count: Counter
	Generic Map ( overflow_count =>7)
	Port Map(
		reset => reset_counter,					-- reset the counter to 0
      counter_clk => clk_in,					-- clock of counter is same as clock of transmitter
      overflow => overflow						-- overflow bit of counter
	);
	
	
	-- process to define the actions in each state
	states:process(clk_in)
	begin
		-- on every rising edge of clock
		if (rising_edge(clk_in)) then
			-- change the present state to old next state
			p_state<=n_state;
			-- depending on the previous next state, (which is now assigned to present state)
			case n_state is
				-- if the state is idle, then high output
				when idle => 
					output <= '1';
					data_sent <= '0';
				
				-- if transmission is to be started, give a low output bit
				when start_transmission =>
					output <= '0';
					data_sent <= '0';
				
				-- after appending 0 bit, start sending data (from output of PISO)
				when data_transmission =>
					output <= out_temp;
					data_sent <= '0';
				
				-- When all the bits are transmitted, give a high output bit
				-- data_sent is made '1' to signify that all bits are transferred
				when stop_transmission =>
					output <= '1';
					data_sent <= '1';
				
			end case;
		end if;
	end process;
	
	-- process to define state transitions
	state_transition: process(send, reset, p_state, overflow)
	begin
		
		-- asynchronus reset which sends the state back to idle
		if (reset='1') then
			n_state <= idle;
		else 
			-- state transitions
			case p_state is 
			
				-- if in idle state, 
				when idle =>
					-- negative edge trigerred send input, which loads input and starts transmission 
					if (send'event and send='0') then 
						n_state <= start_transmission;
						load <='1';
					
					-- else stay in idle state
					else	
						n_state <= idle;

					end if;
					
				-- if transmission is started,
				-- start counting the number of bits outputted, and go to transmission state
				when start_transmission =>
					reset_counter <='1';
					n_state <= data_transmission;
					load <='0';
					
				-- if data is to be transmitted,
				-- count till all the bits are transmitted, and change the state to 'stop_transmission' after 8 bits
				when data_transmission =>
					reset_counter <= '0';
					if (overflow='1') then
						n_state<=stop_transmission;
					else 
						n_state<=data_transmission;
					end if;
				
				-- if all data is transferred, 
				-- go back to idle state
				when stop_transmission =>
					n_state<=idle;
					
				end case;
			end if;
					
	end process;
end Behavioral;

